-- Version: 
-- VHDL Black Box file 
-- 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity MSS_010 is
	generic (
		INIT:std_logic_vector := x"0";
		ACT_UBITS:std_logic_vector := x"0";
		MEMORYFILE:string := "";
		RTC_MAIN_XTL_FREQ:real := 0.0;
		RTC_MAIN_XTL_MODE:string := "";
		DDR_CLK_FREQ:real := 0.0	);
   port( 
       CAN_RXBUS_MGPIO3A_H2F_A : out std_logic;
       CAN_RXBUS_MGPIO3A_H2F_B : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_A : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_B : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_A : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_B : out std_logic;
       CLK_CONFIG_APB : out std_logic;
       COMMS_INT : out std_logic;
       CONFIG_PRESET_N : out std_logic;
       EDAC_ERROR : out std_logic_vector(7 downto 0);
       F_FM0_RDATA : out std_logic_vector(31 downto 0);
       F_FM0_READYOUT : out std_logic;
       F_FM0_RESP : out std_logic;
       F_HM0_ADDR : out std_logic_vector(31 downto 0);
       F_HM0_ENABLE : out std_logic;
       F_HM0_SEL : out std_logic;
       F_HM0_SIZE : out std_logic_vector(1 downto 0);
       F_HM0_TRANS1 : out std_logic;
       F_HM0_WDATA : out std_logic_vector(31 downto 0);
       F_HM0_WRITE : out std_logic;
       FAB_CHRGVBUS : out std_logic;
       FAB_DISCHRGVBUS : out std_logic;
       FAB_DMPULLDOWN : out std_logic;
       FAB_DPPULLDOWN : out std_logic;
       FAB_DRVVBUS : out std_logic;
       FAB_IDPULLUP : out std_logic;
       FAB_OPMODE : out std_logic_vector(1 downto 0);
       FAB_SUSPENDM : out std_logic;
       FAB_TERMSEL : out std_logic;
       FAB_TXVALID : out std_logic;
       FAB_VCONTROL : out std_logic_vector(3 downto 0);
       FAB_VCONTROLLOADM : out std_logic;
       FAB_XCVRSEL : out std_logic_vector(1 downto 0);
       FAB_XDATAOUT : out std_logic_vector(7 downto 0);
       FACC_GLMUX_SEL : out std_logic;
       FIC32_0_MASTER : out std_logic_vector(1 downto 0);
       FIC32_1_MASTER : out std_logic_vector(1 downto 0);
       FPGA_RESET_N : out std_logic;
       GTX_CLK : out std_logic;
       H2F_INTERRUPT : out std_logic_vector(15 downto 0);
       H2F_NMI : out std_logic;
       H2FCALIB : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_A : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_B : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_A : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_B : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_A : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_B : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_A : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_B : out std_logic;
       MDCF : out std_logic;
       MDOENF : out std_logic;
       MDOF : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_A : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_B : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_A : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_B : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_A : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_B : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_A : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_B : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_A : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_B : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_A : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_B : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_A : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_B : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_A : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_B : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_A : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_B : out std_logic;
       MMUART1_DTR_MGPIO12B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_B : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_A : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_B : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_A : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_B : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_A : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_B : out std_logic;
       MPLL_LOCK : out std_logic;
       PER2_FABRIC_PADDR : out std_logic_vector(15 downto 2);
       PER2_FABRIC_PENABLE : out std_logic;
       PER2_FABRIC_PSEL : out std_logic;
       PER2_FABRIC_PWDATA : out std_logic_vector(31 downto 0);
       PER2_FABRIC_PWRITE : out std_logic;
       RTC_MATCH : out std_logic;
       SLEEPDEEP : out std_logic;
       SLEEPHOLDACK : out std_logic;
       SLEEPING : out std_logic;
       SMBALERT_NO0 : out std_logic;
       SMBALERT_NO1 : out std_logic;
       SMBSUS_NO0 : out std_logic;
       SMBSUS_NO1 : out std_logic;
       SPI0_CLK_OUT : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_A : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_B : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_A : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_B : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_A : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_B : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_A : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_B : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_A : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_B : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_A : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_B : out std_logic;
       SPI0_SS4_MGPIO19A_H2F_A : out std_logic;
       SPI0_SS5_MGPIO20A_H2F_A : out std_logic;
       SPI0_SS6_MGPIO21A_H2F_A : out std_logic;
       SPI0_SS7_MGPIO22A_H2F_A : out std_logic;
       SPI1_CLK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_A : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_B : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_A : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_B : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_A : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_B : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_A : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_B : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_A : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_B : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_A : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_B : out std_logic;
       SPI1_SS4_MGPIO17A_H2F_A : out std_logic;
       SPI1_SS5_MGPIO18A_H2F_A : out std_logic;
       SPI1_SS6_MGPIO23A_H2F_A : out std_logic;
       SPI1_SS7_MGPIO24A_H2F_A : out std_logic;
       TCGF : out std_logic_vector(9 downto 0);
       TRACECLK : out std_logic;
       TRACEDATA : out std_logic_vector(3 downto 0);
       TX_CLK : out std_logic;
       TX_ENF : out std_logic;
       TX_ERRF : out std_logic;
       TXCTL_EN_RIF : out std_logic;
       TXD_RIF : out std_logic_vector(3 downto 0);
       TXDF : out std_logic_vector(7 downto 0);
       TXEV : out std_logic;
       WDOGTIMEOUT : out std_logic;
       F_ARREADY_HREADYOUT1 : out std_logic;
       F_AWREADY_HREADYOUT0 : out std_logic;
       F_BID : out std_logic_vector(3 downto 0);
       F_BRESP_HRESP0 : out std_logic_vector(1 downto 0);
       F_BVALID : out std_logic;
       F_RDATA_HRDATA01 : out std_logic_vector(63 downto 0);
       F_RID : out std_logic_vector(3 downto 0);
       F_RLAST : out std_logic;
       F_RRESP_HRESP1 : out std_logic_vector(1 downto 0);
       F_RVALID : out std_logic;
       F_WREADY : out std_logic;
       MDDR_FABRIC_PRDATA : out std_logic_vector(15 downto 0);
       MDDR_FABRIC_PREADY : out std_logic;
       MDDR_FABRIC_PSLVERR : out std_logic;
       CAN_RXBUS_F2H_SCP : in std_logic;
       CAN_TX_EBL_F2H_SCP : in std_logic;
       CAN_TXBUS_F2H_SCP : in std_logic;
       COLF : in std_logic;
       CRSF : in std_logic;
       F2_DMAREADY : in std_logic_vector(1 downto 0);
       F2H_INTERRUPT : in std_logic_vector(15 downto 0);
       F2HCALIB : in std_logic;
       F_DMAREADY : in std_logic_vector(1 downto 0);
       F_FM0_ADDR : in std_logic_vector(31 downto 0);
       F_FM0_ENABLE : in std_logic;
       F_FM0_MASTLOCK : in std_logic;
       F_FM0_READY : in std_logic;
       F_FM0_SEL : in std_logic;
       F_FM0_SIZE : in std_logic_vector(1 downto 0);
       F_FM0_TRANS1 : in std_logic;
       F_FM0_WDATA : in std_logic_vector(31 downto 0);
       F_FM0_WRITE : in std_logic;
       F_HM0_RDATA : in std_logic_vector(31 downto 0);
       F_HM0_READY : in std_logic;
       F_HM0_RESP : in std_logic;
       FAB_AVALID : in std_logic;
       FAB_HOSTDISCON : in std_logic;
       FAB_IDDIG : in std_logic;
       FAB_LINESTATE : in std_logic_vector(1 downto 0);
       FAB_M3_RESET_N : in std_logic;
       FAB_PLL_LOCK : in std_logic;
       FAB_RXACTIVE : in std_logic;
       FAB_RXERROR : in std_logic;
       FAB_RXVALID : in std_logic;
       FAB_RXVALIDH : in std_logic;
       FAB_SESSEND : in std_logic;
       FAB_TXREADY : in std_logic;
       FAB_VBUSVALID : in std_logic;
       FAB_VSTATUS : in std_logic_vector(7 downto 0);
       FAB_XDATAIN : in std_logic_vector(7 downto 0);
       GTX_CLKPF : in std_logic;
       I2C0_BCLK : in std_logic;
       I2C0_SCL_F2H_SCP : in std_logic;
       I2C0_SDA_F2H_SCP : in std_logic;
       I2C1_BCLK : in std_logic;
       I2C1_SCL_F2H_SCP : in std_logic;
       I2C1_SDA_F2H_SCP : in std_logic;
       MDIF : in std_logic;
       MGPIO0A_F2H_GPIN : in std_logic;
       MGPIO10A_F2H_GPIN : in std_logic;
       MGPIO11A_F2H_GPIN : in std_logic;
       MGPIO11B_F2H_GPIN : in std_logic;
       MGPIO12A_F2H_GPIN : in std_logic;
       MGPIO13A_F2H_GPIN : in std_logic;
       MGPIO14A_F2H_GPIN : in std_logic;
       MGPIO15A_F2H_GPIN : in std_logic;
       MGPIO16A_F2H_GPIN : in std_logic;
       MGPIO17B_F2H_GPIN : in std_logic;
       MGPIO18B_F2H_GPIN : in std_logic;
       MGPIO19B_F2H_GPIN : in std_logic;
       MGPIO1A_F2H_GPIN : in std_logic;
       MGPIO20B_F2H_GPIN : in std_logic;
       MGPIO21B_F2H_GPIN : in std_logic;
       MGPIO22B_F2H_GPIN : in std_logic;
       MGPIO24B_F2H_GPIN : in std_logic;
       MGPIO25B_F2H_GPIN : in std_logic;
       MGPIO26B_F2H_GPIN : in std_logic;
       MGPIO27B_F2H_GPIN : in std_logic;
       MGPIO28B_F2H_GPIN : in std_logic;
       MGPIO29B_F2H_GPIN : in std_logic;
       MGPIO2A_F2H_GPIN : in std_logic;
       MGPIO30B_F2H_GPIN : in std_logic;
       MGPIO31B_F2H_GPIN : in std_logic;
       MGPIO3A_F2H_GPIN : in std_logic;
       MGPIO4A_F2H_GPIN : in std_logic;
       MGPIO5A_F2H_GPIN : in std_logic;
       MGPIO6A_F2H_GPIN : in std_logic;
       MGPIO7A_F2H_GPIN : in std_logic;
       MGPIO8A_F2H_GPIN : in std_logic;
       MGPIO9A_F2H_GPIN : in std_logic;
       MMUART0_CTS_F2H_SCP : in std_logic;
       MMUART0_DCD_F2H_SCP : in std_logic;
       MMUART0_DSR_F2H_SCP : in std_logic;
       MMUART0_DTR_F2H_SCP : in std_logic;
       MMUART0_RI_F2H_SCP : in std_logic;
       MMUART0_RTS_F2H_SCP : in std_logic;
       MMUART0_RXD_F2H_SCP : in std_logic;
       MMUART0_SCK_F2H_SCP : in std_logic;
       MMUART0_TXD_F2H_SCP : in std_logic;
       MMUART1_CTS_F2H_SCP : in std_logic;
       MMUART1_DCD_F2H_SCP : in std_logic;
       MMUART1_DSR_F2H_SCP : in std_logic;
       MMUART1_RI_F2H_SCP : in std_logic;
       MMUART1_RTS_F2H_SCP : in std_logic;
       MMUART1_RXD_F2H_SCP : in std_logic;
       MMUART1_SCK_F2H_SCP : in std_logic;
       MMUART1_TXD_F2H_SCP : in std_logic;
       PER2_FABRIC_PRDATA : in std_logic_vector(31 downto 0);
       PER2_FABRIC_PREADY : in std_logic;
       PER2_FABRIC_PSLVERR : in std_logic;
       RCGF : in std_logic_vector(9 downto 0);
       RX_CLKPF : in std_logic;
       RX_DVF : in std_logic;
       RX_ERRF : in std_logic;
       RX_EV : in std_logic;
       RXDF : in std_logic_vector(7 downto 0);
       SLEEPHOLDREQ : in std_logic;
       SMBALERT_NI0 : in std_logic;
       SMBALERT_NI1 : in std_logic;
       SMBSUS_NI0 : in std_logic;
       SMBSUS_NI1 : in std_logic;
       SPI0_CLK_IN : in std_logic;
       SPI0_SDI_F2H_SCP : in std_logic;
       SPI0_SDO_F2H_SCP : in std_logic;
       SPI0_SS0_F2H_SCP : in std_logic;
       SPI0_SS1_F2H_SCP : in std_logic;
       SPI0_SS2_F2H_SCP : in std_logic;
       SPI0_SS3_F2H_SCP : in std_logic;
       SPI1_CLK_IN : in std_logic;
       SPI1_SDI_F2H_SCP : in std_logic;
       SPI1_SDO_F2H_SCP : in std_logic;
       SPI1_SS0_F2H_SCP : in std_logic;
       SPI1_SS1_F2H_SCP : in std_logic;
       SPI1_SS2_F2H_SCP : in std_logic;
       SPI1_SS3_F2H_SCP : in std_logic;
       TX_CLKPF : in std_logic;
       USER_MSS_GPIO_RESET_N : in std_logic;
       USER_MSS_RESET_N : in std_logic;
       XCLK_FAB : in std_logic;
       CLK_BASE : in std_logic;
       CLK_MDDR_APB : in std_logic;
       F_ARADDR_HADDR1 : in std_logic_vector(31 downto 0);
       F_ARBURST_HTRANS1 : in std_logic_vector(1 downto 0);
       F_ARID_HSEL1 : in std_logic_vector(3 downto 0);
       F_ARLEN_HBURST1 : in std_logic_vector(3 downto 0);
       F_ARLOCK_HMASTLOCK1 : in std_logic_vector(1 downto 0);
       F_ARSIZE_HSIZE1 : in std_logic_vector(1 downto 0);
       F_ARVALID_HWRITE1 : in std_logic;
       F_AWADDR_HADDR0 : in std_logic_vector(31 downto 0);
       F_AWBURST_HTRANS0 : in std_logic_vector(1 downto 0);
       F_AWID_HSEL0 : in std_logic_vector(3 downto 0);
       F_AWLEN_HBURST0 : in std_logic_vector(3 downto 0);
       F_AWLOCK_HMASTLOCK0 : in std_logic_vector(1 downto 0);
       F_AWSIZE_HSIZE0 : in std_logic_vector(1 downto 0);
       F_AWVALID_HWRITE0 : in std_logic;
       F_BREADY : in std_logic;
       F_RMW_AXI : in std_logic;
       F_RREADY : in std_logic;
       F_WDATA_HWDATA01 : in std_logic_vector(63 downto 0);
       F_WID_HREADY01 : in std_logic_vector(3 downto 0);
       F_WLAST : in std_logic;
       F_WSTRB : in std_logic_vector(7 downto 0);
       F_WVALID : in std_logic;
       FPGA_MDDR_ARESET_N : in std_logic;
       MDDR_FABRIC_PADDR : in std_logic_vector(10 downto 2);
       MDDR_FABRIC_PENABLE : in std_logic;
       MDDR_FABRIC_PSEL : in std_logic;
       MDDR_FABRIC_PWDATA : in std_logic_vector(15 downto 0);
       MDDR_FABRIC_PWRITE : in std_logic;
       PRESET_N : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN : in std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN : in std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN : in std_logic;
       DM_IN : in std_logic_vector(2 downto 0);
       DRAM_DQ_IN : in std_logic_vector(17 downto 0);
       DRAM_DQS_IN : in std_logic_vector(2 downto 0);
       DRAM_FIFO_WE_IN : in std_logic_vector(1 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN : in std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN : in std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN : in std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN : in std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN : in std_logic;
       MMUART0_DCD_MGPIO22B_IN : in std_logic;
       MMUART0_DSR_MGPIO20B_IN : in std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN : in std_logic;
       MMUART0_RI_MGPIO21B_IN : in std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN : in std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_IN : in std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN : in std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN : in std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN : in std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN : in std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN : in std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN : in std_logic;
       RGMII_MDC_RMII_MDC_IN : in std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN : in std_logic;
       RGMII_RX_CLK_IN : in std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN : in std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN : in std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN : in std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN : in std_logic;
       RGMII_RXD3_USBB_DATA4_IN : in std_logic;
       RGMII_TX_CLK_IN : in std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN : in std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN : in std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN : in std_logic;
       RGMII_TXD2_USBB_DATA5_IN : in std_logic;
       RGMII_TXD3_USBB_DATA6_IN : in std_logic;
       SPI0_SCK_USBA_XCLK_IN : in std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_IN : in std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_IN : in std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_IN : in std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN : in std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN : in std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN : in std_logic;
       SPI1_SCK_IN : in std_logic;
       SPI1_SDI_MGPIO11A_IN : in std_logic;
       SPI1_SDO_MGPIO12A_IN : in std_logic;
       SPI1_SS0_MGPIO13A_IN : in std_logic;
       SPI1_SS1_MGPIO14A_IN : in std_logic;
       SPI1_SS2_MGPIO15A_IN : in std_logic;
       SPI1_SS3_MGPIO16A_IN : in std_logic;
       SPI1_SS4_MGPIO17A_IN : in std_logic;
       SPI1_SS5_MGPIO18A_IN : in std_logic;
       SPI1_SS6_MGPIO23A_IN : in std_logic;
       SPI1_SS7_MGPIO24A_IN : in std_logic;
       USBC_XCLK_IN : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT : out std_logic;
       DRAM_ADDR : out std_logic_vector(15 downto 0);
       DRAM_BA : out std_logic_vector(2 downto 0);
       DRAM_CASN : out std_logic;
       DRAM_CKE : out std_logic;
       DRAM_CLK : out std_logic;
       DRAM_CSN : out std_logic;
       DRAM_DM_RDQS_OUT : out std_logic_vector(2 downto 0);
       DRAM_DQ_OUT : out std_logic_vector(17 downto 0);
       DRAM_DQS_OUT : out std_logic_vector(2 downto 0);
       DRAM_FIFO_WE_OUT : out std_logic_vector(1 downto 0);
       DRAM_ODT : out std_logic;
       DRAM_RASN : out std_logic;
       DRAM_RSTN : out std_logic;
       DRAM_WEN : out std_logic;
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT : out std_logic;
       MMUART0_DCD_MGPIO22B_OUT : out std_logic;
       MMUART0_DSR_MGPIO20B_OUT : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT : out std_logic;
       MMUART0_RI_MGPIO21B_OUT : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT : out std_logic;
       RGMII_MDC_RMII_MDC_OUT : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT : out std_logic;
       RGMII_RX_CLK_OUT : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT : out std_logic;
       RGMII_RXD3_USBB_DATA4_OUT : out std_logic;
       RGMII_TX_CLK_OUT : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT : out std_logic;
       RGMII_TXD2_USBB_DATA5_OUT : out std_logic;
       RGMII_TXD3_USBB_DATA6_OUT : out std_logic;
       SPI0_SCK_USBA_XCLK_OUT : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OUT : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT : out std_logic;
       SPI1_SCK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_OUT : out std_logic;
       SPI1_SDO_MGPIO12A_OUT : out std_logic;
       SPI1_SS0_MGPIO13A_OUT : out std_logic;
       SPI1_SS1_MGPIO14A_OUT : out std_logic;
       SPI1_SS2_MGPIO15A_OUT : out std_logic;
       SPI1_SS3_MGPIO16A_OUT : out std_logic;
       SPI1_SS4_MGPIO17A_OUT : out std_logic;
       SPI1_SS5_MGPIO18A_OUT : out std_logic;
       SPI1_SS6_MGPIO23A_OUT : out std_logic;
       SPI1_SS7_MGPIO24A_OUT : out std_logic;
       USBC_XCLK_OUT : out std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE : out std_logic;
       DM_OE : out std_logic_vector(2 downto 0);
       DRAM_DQ_OE : out std_logic_vector(17 downto 0);
       DRAM_DQS_OE : out std_logic_vector(2 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE : out std_logic;
       MMUART0_DCD_MGPIO22B_OE : out std_logic;
       MMUART0_DSR_MGPIO20B_OE : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE : out std_logic;
       MMUART0_RI_MGPIO21B_OE : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OE : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE : out std_logic;
       RGMII_MDC_RMII_MDC_OE : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE : out std_logic;
       RGMII_RX_CLK_OE : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE : out std_logic;
       RGMII_RXD3_USBB_DATA4_OE : out std_logic;
       RGMII_TX_CLK_OE : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE : out std_logic;
       RGMII_TXD2_USBB_DATA5_OE : out std_logic;
       RGMII_TXD3_USBB_DATA6_OE : out std_logic;
       SPI0_SCK_USBA_XCLK_OE : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OE : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OE : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OE : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE : out std_logic;
       SPI1_SCK_OE : out std_logic;
       SPI1_SDI_MGPIO11A_OE : out std_logic;
       SPI1_SDO_MGPIO12A_OE : out std_logic;
       SPI1_SS0_MGPIO13A_OE : out std_logic;
       SPI1_SS1_MGPIO14A_OE : out std_logic;
       SPI1_SS2_MGPIO15A_OE : out std_logic;
       SPI1_SS3_MGPIO16A_OE : out std_logic;
       SPI1_SS4_MGPIO17A_OE : out std_logic;
       SPI1_SS5_MGPIO18A_OE : out std_logic;
       SPI1_SS6_MGPIO23A_OE : out std_logic;
       SPI1_SS7_MGPIO24A_OE : out std_logic;
       USBC_XCLK_OE : out std_logic
   );
end MSS_010;
architecture DEF_ARCH of MSS_010 is 

   attribute syn_black_box : boolean;
   attribute syn_black_box of DEF_ARCH : architecture is true;
   attribute syn_tsu0: string;
   attribute syn_tsu0 of DEF_ARCH : architecture is " CAN_RXBUS_F2H_SCP->CLK_BASE = 1.047";
   attribute syn_tsu1: string;
   attribute syn_tsu1 of DEF_ARCH : architecture is " F2HCALIB->CLK_BASE = 0.39";
   attribute syn_tsu2: string;
   attribute syn_tsu2 of DEF_ARCH : architecture is " F2H_INTERRUPT[0]->CLK_BASE = 0.858";
   attribute syn_tsu3: string;
   attribute syn_tsu3 of DEF_ARCH : architecture is " F2H_INTERRUPT[10]->CLK_BASE = 1.07";
   attribute syn_tsu4: string;
   attribute syn_tsu4 of DEF_ARCH : architecture is " F2H_INTERRUPT[11]->CLK_BASE = 1.049";
   attribute syn_tsu5: string;
   attribute syn_tsu5 of DEF_ARCH : architecture is " F2H_INTERRUPT[12]->CLK_BASE = 0.967";
   attribute syn_tsu6: string;
   attribute syn_tsu6 of DEF_ARCH : architecture is " F2H_INTERRUPT[13]->CLK_BASE = 1.024";
   attribute syn_tsu7: string;
   attribute syn_tsu7 of DEF_ARCH : architecture is " F2H_INTERRUPT[14]->CLK_BASE = 1.077";
   attribute syn_tsu8: string;
   attribute syn_tsu8 of DEF_ARCH : architecture is " F2H_INTERRUPT[15]->CLK_BASE = 0.989";
   attribute syn_tsu9: string;
   attribute syn_tsu9 of DEF_ARCH : architecture is " F2H_INTERRUPT[1]->CLK_BASE = 0.824";
   attribute syn_tsu10: string;
   attribute syn_tsu10 of DEF_ARCH : architecture is " F2H_INTERRUPT[2]->CLK_BASE = 0.791";
   attribute syn_tsu11: string;
   attribute syn_tsu11 of DEF_ARCH : architecture is " F2H_INTERRUPT[3]->CLK_BASE = 0.907";
   attribute syn_tsu12: string;
   attribute syn_tsu12 of DEF_ARCH : architecture is " F2H_INTERRUPT[4]->CLK_BASE = 0.803";
   attribute syn_tsu13: string;
   attribute syn_tsu13 of DEF_ARCH : architecture is " F2H_INTERRUPT[5]->CLK_BASE = 0.911";
   attribute syn_tsu14: string;
   attribute syn_tsu14 of DEF_ARCH : architecture is " F2H_INTERRUPT[6]->CLK_BASE = 0.864";
   attribute syn_tsu15: string;
   attribute syn_tsu15 of DEF_ARCH : architecture is " F2H_INTERRUPT[7]->CLK_BASE = 0.902";
   attribute syn_tsu16: string;
   attribute syn_tsu16 of DEF_ARCH : architecture is " F2H_INTERRUPT[8]->CLK_BASE = 0.882";
   attribute syn_tsu17: string;
   attribute syn_tsu17 of DEF_ARCH : architecture is " F2H_INTERRUPT[9]->CLK_BASE = 0.825";
   attribute syn_tsu18: string;
   attribute syn_tsu18 of DEF_ARCH : architecture is " F_FM0_ADDR[0]->CLK_BASE = 0.915";
   attribute syn_tsu19: string;
   attribute syn_tsu19 of DEF_ARCH : architecture is " F_FM0_ADDR[10]->CLK_BASE = 0.848";
   attribute syn_tsu20: string;
   attribute syn_tsu20 of DEF_ARCH : architecture is " F_FM0_ADDR[11]->CLK_BASE = 0.957";
   attribute syn_tsu21: string;
   attribute syn_tsu21 of DEF_ARCH : architecture is " F_FM0_ADDR[12]->CLK_BASE = 0.967";
   attribute syn_tsu22: string;
   attribute syn_tsu22 of DEF_ARCH : architecture is " F_FM0_ADDR[13]->CLK_BASE = 1.194";
   attribute syn_tsu23: string;
   attribute syn_tsu23 of DEF_ARCH : architecture is " F_FM0_ADDR[14]->CLK_BASE = 1.105";
   attribute syn_tsu24: string;
   attribute syn_tsu24 of DEF_ARCH : architecture is " F_FM0_ADDR[15]->CLK_BASE = 1.093";
   attribute syn_tsu25: string;
   attribute syn_tsu25 of DEF_ARCH : architecture is " F_FM0_ADDR[16]->CLK_BASE = 1.071";
   attribute syn_tsu26: string;
   attribute syn_tsu26 of DEF_ARCH : architecture is " F_FM0_ADDR[17]->CLK_BASE = 1.001";
   attribute syn_tsu27: string;
   attribute syn_tsu27 of DEF_ARCH : architecture is " F_FM0_ADDR[18]->CLK_BASE = 1.068";
   attribute syn_tsu28: string;
   attribute syn_tsu28 of DEF_ARCH : architecture is " F_FM0_ADDR[19]->CLK_BASE = 0.571";
   attribute syn_tsu29: string;
   attribute syn_tsu29 of DEF_ARCH : architecture is " F_FM0_ADDR[1]->CLK_BASE = 0.801";
   attribute syn_tsu30: string;
   attribute syn_tsu30 of DEF_ARCH : architecture is " F_FM0_ADDR[20]->CLK_BASE = 0.879";
   attribute syn_tsu31: string;
   attribute syn_tsu31 of DEF_ARCH : architecture is " F_FM0_ADDR[21]->CLK_BASE = 0.532";
   attribute syn_tsu32: string;
   attribute syn_tsu32 of DEF_ARCH : architecture is " F_FM0_ADDR[22]->CLK_BASE = 0.878";
   attribute syn_tsu33: string;
   attribute syn_tsu33 of DEF_ARCH : architecture is " F_FM0_ADDR[23]->CLK_BASE = 0.575";
   attribute syn_tsu34: string;
   attribute syn_tsu34 of DEF_ARCH : architecture is " F_FM0_ADDR[24]->CLK_BASE = 0.596";
   attribute syn_tsu35: string;
   attribute syn_tsu35 of DEF_ARCH : architecture is " F_FM0_ADDR[25]->CLK_BASE = 0.663";
   attribute syn_tsu36: string;
   attribute syn_tsu36 of DEF_ARCH : architecture is " F_FM0_ADDR[26]->CLK_BASE = 0.712";
   attribute syn_tsu37: string;
   attribute syn_tsu37 of DEF_ARCH : architecture is " F_FM0_ADDR[27]->CLK_BASE = 1.073";
   attribute syn_tsu38: string;
   attribute syn_tsu38 of DEF_ARCH : architecture is " F_FM0_ADDR[28]->CLK_BASE = 0.696";
   attribute syn_tsu39: string;
   attribute syn_tsu39 of DEF_ARCH : architecture is " F_FM0_ADDR[29]->CLK_BASE = 0.399";
   attribute syn_tsu40: string;
   attribute syn_tsu40 of DEF_ARCH : architecture is " F_FM0_ADDR[2]->CLK_BASE = 0.331";
   attribute syn_tsu41: string;
   attribute syn_tsu41 of DEF_ARCH : architecture is " F_FM0_ADDR[30]->CLK_BASE = 0.582";
   attribute syn_tsu42: string;
   attribute syn_tsu42 of DEF_ARCH : architecture is " F_FM0_ADDR[31]->CLK_BASE = 0.479";
   attribute syn_tsu43: string;
   attribute syn_tsu43 of DEF_ARCH : architecture is " F_FM0_ADDR[3]->CLK_BASE = 0.956";
   attribute syn_tsu44: string;
   attribute syn_tsu44 of DEF_ARCH : architecture is " F_FM0_ADDR[4]->CLK_BASE = 1.273";
   attribute syn_tsu45: string;
   attribute syn_tsu45 of DEF_ARCH : architecture is " F_FM0_ADDR[5]->CLK_BASE = 0.844";
   attribute syn_tsu46: string;
   attribute syn_tsu46 of DEF_ARCH : architecture is " F_FM0_ADDR[6]->CLK_BASE = 1.139";
   attribute syn_tsu47: string;
   attribute syn_tsu47 of DEF_ARCH : architecture is " F_FM0_ADDR[7]->CLK_BASE = 1.031";
   attribute syn_tsu48: string;
   attribute syn_tsu48 of DEF_ARCH : architecture is " F_FM0_ADDR[8]->CLK_BASE = 1.018";
   attribute syn_tsu49: string;
   attribute syn_tsu49 of DEF_ARCH : architecture is " F_FM0_ADDR[9]->CLK_BASE = 0.786";
   attribute syn_tsu50: string;
   attribute syn_tsu50 of DEF_ARCH : architecture is " F_FM0_ENABLE->CLK_BASE = 1.163";
   attribute syn_tsu51: string;
   attribute syn_tsu51 of DEF_ARCH : architecture is " F_FM0_SEL->CLK_BASE = 1.409";
   attribute syn_tsu52: string;
   attribute syn_tsu52 of DEF_ARCH : architecture is " F_FM0_WDATA[0]->CLK_BASE = 0.131";
   attribute syn_tsu53: string;
   attribute syn_tsu53 of DEF_ARCH : architecture is " F_FM0_WDATA[10]->CLK_BASE = 0.158";
   attribute syn_tsu54: string;
   attribute syn_tsu54 of DEF_ARCH : architecture is " F_FM0_WDATA[11]->CLK_BASE = 0.086";
   attribute syn_tsu55: string;
   attribute syn_tsu55 of DEF_ARCH : architecture is " F_FM0_WDATA[12]->CLK_BASE = 0.098";
   attribute syn_tsu56: string;
   attribute syn_tsu56 of DEF_ARCH : architecture is " F_FM0_WDATA[13]->CLK_BASE = 0.093";
   attribute syn_tsu57: string;
   attribute syn_tsu57 of DEF_ARCH : architecture is " F_FM0_WDATA[14]->CLK_BASE = 0.14";
   attribute syn_tsu58: string;
   attribute syn_tsu58 of DEF_ARCH : architecture is " F_FM0_WDATA[15]->CLK_BASE = 0.126";
   attribute syn_tsu59: string;
   attribute syn_tsu59 of DEF_ARCH : architecture is " F_FM0_WDATA[16]->CLK_BASE = 0.103";
   attribute syn_tsu60: string;
   attribute syn_tsu60 of DEF_ARCH : architecture is " F_FM0_WDATA[17]->CLK_BASE = 0.107";
   attribute syn_tsu61: string;
   attribute syn_tsu61 of DEF_ARCH : architecture is " F_FM0_WDATA[18]->CLK_BASE = 0.152";
   attribute syn_tsu62: string;
   attribute syn_tsu62 of DEF_ARCH : architecture is " F_FM0_WDATA[19]->CLK_BASE = 0.13";
   attribute syn_tsu63: string;
   attribute syn_tsu63 of DEF_ARCH : architecture is " F_FM0_WDATA[1]->CLK_BASE = 0.087";
   attribute syn_tsu64: string;
   attribute syn_tsu64 of DEF_ARCH : architecture is " F_FM0_WDATA[20]->CLK_BASE = 0.108";
   attribute syn_tsu65: string;
   attribute syn_tsu65 of DEF_ARCH : architecture is " F_FM0_WDATA[21]->CLK_BASE = 0.054";
   attribute syn_tsu66: string;
   attribute syn_tsu66 of DEF_ARCH : architecture is " F_FM0_WDATA[22]->CLK_BASE = 0.052";
   attribute syn_tsu67: string;
   attribute syn_tsu67 of DEF_ARCH : architecture is " F_FM0_WDATA[23]->CLK_BASE = 0.084";
   attribute syn_tsu68: string;
   attribute syn_tsu68 of DEF_ARCH : architecture is " F_FM0_WDATA[24]->CLK_BASE = 0.094";
   attribute syn_tsu69: string;
   attribute syn_tsu69 of DEF_ARCH : architecture is " F_FM0_WDATA[25]->CLK_BASE = 0.177";
   attribute syn_tsu70: string;
   attribute syn_tsu70 of DEF_ARCH : architecture is " F_FM0_WDATA[26]->CLK_BASE = 0.117";
   attribute syn_tsu71: string;
   attribute syn_tsu71 of DEF_ARCH : architecture is " F_FM0_WDATA[27]->CLK_BASE = 0.096";
   attribute syn_tsu72: string;
   attribute syn_tsu72 of DEF_ARCH : architecture is " F_FM0_WDATA[28]->CLK_BASE = 0.157";
   attribute syn_tsu73: string;
   attribute syn_tsu73 of DEF_ARCH : architecture is " F_FM0_WDATA[29]->CLK_BASE = 0.115";
   attribute syn_tsu74: string;
   attribute syn_tsu74 of DEF_ARCH : architecture is " F_FM0_WDATA[2]->CLK_BASE = 0.059";
   attribute syn_tsu75: string;
   attribute syn_tsu75 of DEF_ARCH : architecture is " F_FM0_WDATA[30]->CLK_BASE = 0.081";
   attribute syn_tsu76: string;
   attribute syn_tsu76 of DEF_ARCH : architecture is " F_FM0_WDATA[31]->CLK_BASE = 0.126";
   attribute syn_tsu77: string;
   attribute syn_tsu77 of DEF_ARCH : architecture is " F_FM0_WDATA[3]->CLK_BASE = 0.096";
   attribute syn_tsu78: string;
   attribute syn_tsu78 of DEF_ARCH : architecture is " F_FM0_WDATA[4]->CLK_BASE = 0.055";
   attribute syn_tsu79: string;
   attribute syn_tsu79 of DEF_ARCH : architecture is " F_FM0_WDATA[5]->CLK_BASE = 0.115";
   attribute syn_tsu80: string;
   attribute syn_tsu80 of DEF_ARCH : architecture is " F_FM0_WDATA[6]->CLK_BASE = 0.082";
   attribute syn_tsu81: string;
   attribute syn_tsu81 of DEF_ARCH : architecture is " F_FM0_WDATA[7]->CLK_BASE = 0.125";
   attribute syn_tsu82: string;
   attribute syn_tsu82 of DEF_ARCH : architecture is " F_FM0_WDATA[8]->CLK_BASE = 0.121";
   attribute syn_tsu83: string;
   attribute syn_tsu83 of DEF_ARCH : architecture is " F_FM0_WDATA[9]->CLK_BASE = 0.074";
   attribute syn_tsu84: string;
   attribute syn_tsu84 of DEF_ARCH : architecture is " F_FM0_WRITE->CLK_BASE = 0.967";
   attribute syn_tsu85: string;
   attribute syn_tsu85 of DEF_ARCH : architecture is " F_HM0_RDATA[0]->CLK_BASE = 0.367";
   attribute syn_tsu86: string;
   attribute syn_tsu86 of DEF_ARCH : architecture is " F_HM0_RDATA[10]->CLK_BASE = 0.244";
   attribute syn_tsu87: string;
   attribute syn_tsu87 of DEF_ARCH : architecture is " F_HM0_RDATA[11]->CLK_BASE = 0.329";
   attribute syn_tsu88: string;
   attribute syn_tsu88 of DEF_ARCH : architecture is " F_HM0_RDATA[12]->CLK_BASE = 0.273";
   attribute syn_tsu89: string;
   attribute syn_tsu89 of DEF_ARCH : architecture is " F_HM0_RDATA[13]->CLK_BASE = 0.341";
   attribute syn_tsu90: string;
   attribute syn_tsu90 of DEF_ARCH : architecture is " F_HM0_RDATA[14]->CLK_BASE = 0.285";
   attribute syn_tsu91: string;
   attribute syn_tsu91 of DEF_ARCH : architecture is " F_HM0_RDATA[15]->CLK_BASE = 0.276";
   attribute syn_tsu92: string;
   attribute syn_tsu92 of DEF_ARCH : architecture is " F_HM0_RDATA[16]->CLK_BASE = 0.333";
   attribute syn_tsu93: string;
   attribute syn_tsu93 of DEF_ARCH : architecture is " F_HM0_RDATA[17]->CLK_BASE = 0.3";
   attribute syn_tsu94: string;
   attribute syn_tsu94 of DEF_ARCH : architecture is " F_HM0_RDATA[18]->CLK_BASE = 0.227";
   attribute syn_tsu95: string;
   attribute syn_tsu95 of DEF_ARCH : architecture is " F_HM0_RDATA[19]->CLK_BASE = 0.284";
   attribute syn_tsu96: string;
   attribute syn_tsu96 of DEF_ARCH : architecture is " F_HM0_RDATA[1]->CLK_BASE = 0.289";
   attribute syn_tsu97: string;
   attribute syn_tsu97 of DEF_ARCH : architecture is " F_HM0_RDATA[20]->CLK_BASE = 0.297";
   attribute syn_tsu98: string;
   attribute syn_tsu98 of DEF_ARCH : architecture is " F_HM0_RDATA[21]->CLK_BASE = 0.321";
   attribute syn_tsu99: string;
   attribute syn_tsu99 of DEF_ARCH : architecture is " F_HM0_RDATA[22]->CLK_BASE = 0.327";
   attribute syn_tsu100: string;
   attribute syn_tsu100 of DEF_ARCH : architecture is " F_HM0_RDATA[23]->CLK_BASE = 0.384";
   attribute syn_tsu101: string;
   attribute syn_tsu101 of DEF_ARCH : architecture is " F_HM0_RDATA[24]->CLK_BASE = 0.296";
   attribute syn_tsu102: string;
   attribute syn_tsu102 of DEF_ARCH : architecture is " F_HM0_RDATA[25]->CLK_BASE = 0.264";
   attribute syn_tsu103: string;
   attribute syn_tsu103 of DEF_ARCH : architecture is " F_HM0_RDATA[26]->CLK_BASE = 0.22";
   attribute syn_tsu104: string;
   attribute syn_tsu104 of DEF_ARCH : architecture is " F_HM0_RDATA[27]->CLK_BASE = 0.278";
   attribute syn_tsu105: string;
   attribute syn_tsu105 of DEF_ARCH : architecture is " F_HM0_RDATA[28]->CLK_BASE = 0.285";
   attribute syn_tsu106: string;
   attribute syn_tsu106 of DEF_ARCH : architecture is " F_HM0_RDATA[29]->CLK_BASE = 0.358";
   attribute syn_tsu107: string;
   attribute syn_tsu107 of DEF_ARCH : architecture is " F_HM0_RDATA[2]->CLK_BASE = 0.263";
   attribute syn_tsu108: string;
   attribute syn_tsu108 of DEF_ARCH : architecture is " F_HM0_RDATA[30]->CLK_BASE = 0.354";
   attribute syn_tsu109: string;
   attribute syn_tsu109 of DEF_ARCH : architecture is " F_HM0_RDATA[31]->CLK_BASE = 0.252";
   attribute syn_tsu110: string;
   attribute syn_tsu110 of DEF_ARCH : architecture is " F_HM0_RDATA[3]->CLK_BASE = 0.525";
   attribute syn_tsu111: string;
   attribute syn_tsu111 of DEF_ARCH : architecture is " F_HM0_RDATA[4]->CLK_BASE = 0.459";
   attribute syn_tsu112: string;
   attribute syn_tsu112 of DEF_ARCH : architecture is " F_HM0_RDATA[5]->CLK_BASE = 0.303";
   attribute syn_tsu113: string;
   attribute syn_tsu113 of DEF_ARCH : architecture is " F_HM0_RDATA[6]->CLK_BASE = 0.328";
   attribute syn_tsu114: string;
   attribute syn_tsu114 of DEF_ARCH : architecture is " F_HM0_RDATA[7]->CLK_BASE = 0.196";
   attribute syn_tsu115: string;
   attribute syn_tsu115 of DEF_ARCH : architecture is " F_HM0_RDATA[8]->CLK_BASE = 0.308";
   attribute syn_tsu116: string;
   attribute syn_tsu116 of DEF_ARCH : architecture is " F_HM0_RDATA[9]->CLK_BASE = 0.396";
   attribute syn_tsu117: string;
   attribute syn_tsu117 of DEF_ARCH : architecture is " F_HM0_READY->CLK_BASE = 1.514";
   attribute syn_tsu118: string;
   attribute syn_tsu118 of DEF_ARCH : architecture is " F_HM0_RESP->CLK_BASE = 0.921";
   attribute syn_tsu119: string;
   attribute syn_tsu119 of DEF_ARCH : architecture is " I2C0_SDA_F2H_SCP->I2C0_SCL_F2H_SCP = 0.214";
   attribute syn_tsu120: string;
   attribute syn_tsu120 of DEF_ARCH : architecture is " I2C1_SDA_F2H_SCP->I2C1_SCL_F2H_SCP = 0.23";
   attribute syn_tsu121: string;
   attribute syn_tsu121 of DEF_ARCH : architecture is " MGPIO0A_F2H_GPIN->CLK_BASE = 0.881";
   attribute syn_tsu122: string;
   attribute syn_tsu122 of DEF_ARCH : architecture is " MGPIO10A_F2H_GPIN->CLK_BASE = 1.068";
   attribute syn_tsu123: string;
   attribute syn_tsu123 of DEF_ARCH : architecture is " MGPIO11A_F2H_GPIN->CLK_BASE = 0.325";
   attribute syn_tsu124: string;
   attribute syn_tsu124 of DEF_ARCH : architecture is " MGPIO11B_F2H_GPIN->CLK_BASE = 0.381";
   attribute syn_tsu125: string;
   attribute syn_tsu125 of DEF_ARCH : architecture is " MGPIO12A_F2H_GPIN->CLK_BASE = 0.385";
   attribute syn_tsu126: string;
   attribute syn_tsu126 of DEF_ARCH : architecture is " MGPIO13A_F2H_GPIN->CLK_BASE = 0.463";
   attribute syn_tsu127: string;
   attribute syn_tsu127 of DEF_ARCH : architecture is " MGPIO14A_F2H_GPIN->CLK_BASE = 0.379";
   attribute syn_tsu128: string;
   attribute syn_tsu128 of DEF_ARCH : architecture is " MGPIO15A_F2H_GPIN->CLK_BASE = 0.414";
   attribute syn_tsu129: string;
   attribute syn_tsu129 of DEF_ARCH : architecture is " MGPIO16A_F2H_GPIN->CLK_BASE = 0.358";
   attribute syn_tsu130: string;
   attribute syn_tsu130 of DEF_ARCH : architecture is " MGPIO17B_F2H_GPIN->CLK_BASE = 0.477";
   attribute syn_tsu131: string;
   attribute syn_tsu131 of DEF_ARCH : architecture is " MGPIO18B_F2H_GPIN->CLK_BASE = 0.5";
   attribute syn_tsu132: string;
   attribute syn_tsu132 of DEF_ARCH : architecture is " MGPIO19B_F2H_GPIN->CLK_BASE = 0.521";
   attribute syn_tsu133: string;
   attribute syn_tsu133 of DEF_ARCH : architecture is " MGPIO1A_F2H_GPIN->CLK_BASE = 0.435";
   attribute syn_tsu134: string;
   attribute syn_tsu134 of DEF_ARCH : architecture is " MGPIO20B_F2H_GPIN->CLK_BASE = 0.468";
   attribute syn_tsu135: string;
   attribute syn_tsu135 of DEF_ARCH : architecture is " MGPIO21B_F2H_GPIN->CLK_BASE = 0.507";
   attribute syn_tsu136: string;
   attribute syn_tsu136 of DEF_ARCH : architecture is " MGPIO22B_F2H_GPIN->CLK_BASE = 0.473";
   attribute syn_tsu137: string;
   attribute syn_tsu137 of DEF_ARCH : architecture is " MGPIO24B_F2H_GPIN->CLK_BASE = 0.381";
   attribute syn_tsu138: string;
   attribute syn_tsu138 of DEF_ARCH : architecture is " MGPIO25B_F2H_GPIN->CLK_BASE = 0.787";
   attribute syn_tsu139: string;
   attribute syn_tsu139 of DEF_ARCH : architecture is " MGPIO26B_F2H_GPIN->CLK_BASE = 0.727";
   attribute syn_tsu140: string;
   attribute syn_tsu140 of DEF_ARCH : architecture is " MGPIO27B_F2H_GPIN->CLK_BASE = 1.08";
   attribute syn_tsu141: string;
   attribute syn_tsu141 of DEF_ARCH : architecture is " MGPIO28B_F2H_GPIN->CLK_BASE = 1.311";
   attribute syn_tsu142: string;
   attribute syn_tsu142 of DEF_ARCH : architecture is " MGPIO29B_F2H_GPIN->CLK_BASE = 1.047";
   attribute syn_tsu143: string;
   attribute syn_tsu143 of DEF_ARCH : architecture is " MGPIO2A_F2H_GPIN->CLK_BASE = 0.746";
   attribute syn_tsu144: string;
   attribute syn_tsu144 of DEF_ARCH : architecture is " MGPIO30B_F2H_GPIN->CLK_BASE = 0.888";
   attribute syn_tsu145: string;
   attribute syn_tsu145 of DEF_ARCH : architecture is " MGPIO31B_F2H_GPIN->CLK_BASE = 0.895";
   attribute syn_tsu146: string;
   attribute syn_tsu146 of DEF_ARCH : architecture is " MGPIO3A_F2H_GPIN->CLK_BASE = 1.046";
   attribute syn_tsu147: string;
   attribute syn_tsu147 of DEF_ARCH : architecture is " MGPIO4A_F2H_GPIN->CLK_BASE = 0.886";
   attribute syn_tsu148: string;
   attribute syn_tsu148 of DEF_ARCH : architecture is " MGPIO5A_F2H_GPIN->CLK_BASE = 0.654";
   attribute syn_tsu149: string;
   attribute syn_tsu149 of DEF_ARCH : architecture is " MGPIO6A_F2H_GPIN->CLK_BASE = 0.704";
   attribute syn_tsu150: string;
   attribute syn_tsu150 of DEF_ARCH : architecture is " MGPIO7A_F2H_GPIN->CLK_BASE = 0.759";
   attribute syn_tsu151: string;
   attribute syn_tsu151 of DEF_ARCH : architecture is " MGPIO8A_F2H_GPIN->CLK_BASE = 0.769";
   attribute syn_tsu152: string;
   attribute syn_tsu152 of DEF_ARCH : architecture is " MGPIO9A_F2H_GPIN->CLK_BASE = 0.68";
   attribute syn_tsu153: string;
   attribute syn_tsu153 of DEF_ARCH : architecture is " MMUART0_CTS_F2H_SCP->CLK_BASE = 0.629";
   attribute syn_tsu154: string;
   attribute syn_tsu154 of DEF_ARCH : architecture is " MMUART0_DCD_F2H_SCP->CLK_BASE = 0.655";
   attribute syn_tsu155: string;
   attribute syn_tsu155 of DEF_ARCH : architecture is " MMUART0_DSR_F2H_SCP->CLK_BASE = 0.781";
   attribute syn_tsu156: string;
   attribute syn_tsu156 of DEF_ARCH : architecture is " MMUART0_RI_F2H_SCP->CLK_BASE = 0.486";
   attribute syn_tsu157: string;
   attribute syn_tsu157 of DEF_ARCH : architecture is " MMUART0_RXD_F2H_SCP->CLK_BASE = 0.559";
   attribute syn_tsu158: string;
   attribute syn_tsu158 of DEF_ARCH : architecture is " MMUART0_SCK_F2H_SCP->CLK_BASE = 0.653";
   attribute syn_tsu159: string;
   attribute syn_tsu159 of DEF_ARCH : architecture is " MMUART0_TXD_F2H_SCP->CLK_BASE = 0.608";
   attribute syn_tsu160: string;
   attribute syn_tsu160 of DEF_ARCH : architecture is " MMUART1_CTS_F2H_SCP->CLK_BASE = 0.956";
   attribute syn_tsu161: string;
   attribute syn_tsu161 of DEF_ARCH : architecture is " MMUART1_DCD_F2H_SCP->CLK_BASE = 1.076";
   attribute syn_tsu162: string;
   attribute syn_tsu162 of DEF_ARCH : architecture is " MMUART1_DSR_F2H_SCP->CLK_BASE = 1.014";
   attribute syn_tsu163: string;
   attribute syn_tsu163 of DEF_ARCH : architecture is " MMUART1_RI_F2H_SCP->CLK_BASE = 0.66";
   attribute syn_tsu164: string;
   attribute syn_tsu164 of DEF_ARCH : architecture is " MMUART1_RXD_F2H_SCP->CLK_BASE = 0.661";
   attribute syn_tsu165: string;
   attribute syn_tsu165 of DEF_ARCH : architecture is " MMUART1_SCK_F2H_SCP->CLK_BASE = 1.057";
   attribute syn_tsu166: string;
   attribute syn_tsu166 of DEF_ARCH : architecture is " MMUART1_TXD_F2H_SCP->CLK_BASE = 0.649";
   attribute syn_tsu167: string;
   attribute syn_tsu167 of DEF_ARCH : architecture is " SMBALERT_NI0->I2C0_SCL_F2H_SCP = 0";
   attribute syn_tsu168: string;
   attribute syn_tsu168 of DEF_ARCH : architecture is " SMBALERT_NI1->I2C1_SCL_F2H_SCP = 0";
   attribute syn_tsu169: string;
   attribute syn_tsu169 of DEF_ARCH : architecture is " SMBSUS_NI0->I2C0_SCL_F2H_SCP = 0";
   attribute syn_tsu170: string;
   attribute syn_tsu170 of DEF_ARCH : architecture is " SMBSUS_NI1->I2C1_SCL_F2H_SCP = 0";
   attribute syn_tsu171: string;
   attribute syn_tsu171 of DEF_ARCH : architecture is " SPI0_SDI_F2H_SCP->SPI0_CLK_IN = 1.304";
   attribute syn_tsu172: string;
   attribute syn_tsu172 of DEF_ARCH : architecture is " SPI1_SDI_F2H_SCP->SPI1_CLK_IN = 1.418";
   attribute syn_tco0: string;
   attribute syn_tco0 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_A = 3.276";
   attribute syn_tco1: string;
   attribute syn_tco1 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_B = 3.202";
   attribute syn_tco2: string;
   attribute syn_tco2 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_A = 3.179";
   attribute syn_tco3: string;
   attribute syn_tco3 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_B = 3.083";
   attribute syn_tco4: string;
   attribute syn_tco4 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT = 4.272";
   attribute syn_tco5: string;
   attribute syn_tco5 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_A = 3.308";
   attribute syn_tco6: string;
   attribute syn_tco6 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_B = 3.278";
   attribute syn_tco7: string;
   attribute syn_tco7 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT = 3.933";
   attribute syn_tco8: string;
   attribute syn_tco8 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[0] = 3.860";
   attribute syn_tco9: string;
   attribute syn_tco9 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[10] = 3.888";
   attribute syn_tco10: string;
   attribute syn_tco10 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[11] = 4.003";
   attribute syn_tco11: string;
   attribute syn_tco11 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[12] = 3.918";
   attribute syn_tco12: string;
   attribute syn_tco12 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[13] = 3.880";
   attribute syn_tco13: string;
   attribute syn_tco13 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[14] = 3.880";
   attribute syn_tco14: string;
   attribute syn_tco14 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[15] = 3.874";
   attribute syn_tco15: string;
   attribute syn_tco15 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[16] = 3.907";
   attribute syn_tco16: string;
   attribute syn_tco16 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[17] = 4.105";
   attribute syn_tco17: string;
   attribute syn_tco17 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[18] = 3.871";
   attribute syn_tco18: string;
   attribute syn_tco18 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[19] = 4.023";
   attribute syn_tco19: string;
   attribute syn_tco19 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[1] = 3.940";
   attribute syn_tco20: string;
   attribute syn_tco20 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[20] = 3.776";
   attribute syn_tco21: string;
   attribute syn_tco21 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[21] = 3.731";
   attribute syn_tco22: string;
   attribute syn_tco22 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[22] = 3.762";
   attribute syn_tco23: string;
   attribute syn_tco23 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[23] = 3.763";
   attribute syn_tco24: string;
   attribute syn_tco24 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[24] = 3.784";
   attribute syn_tco25: string;
   attribute syn_tco25 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[25] = 3.780";
   attribute syn_tco26: string;
   attribute syn_tco26 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[26] = 3.885";
   attribute syn_tco27: string;
   attribute syn_tco27 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[27] = 3.778";
   attribute syn_tco28: string;
   attribute syn_tco28 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[28] = 3.769";
   attribute syn_tco29: string;
   attribute syn_tco29 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[29] = 3.761";
   attribute syn_tco30: string;
   attribute syn_tco30 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[2] = 3.907";
   attribute syn_tco31: string;
   attribute syn_tco31 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[30] = 4.038";
   attribute syn_tco32: string;
   attribute syn_tco32 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[31] = 3.902";
   attribute syn_tco33: string;
   attribute syn_tco33 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[3] = 3.949";
   attribute syn_tco34: string;
   attribute syn_tco34 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[4] = 3.956";
   attribute syn_tco35: string;
   attribute syn_tco35 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[5] = 4.077";
   attribute syn_tco36: string;
   attribute syn_tco36 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[6] = 3.939";
   attribute syn_tco37: string;
   attribute syn_tco37 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[7] = 3.924";
   attribute syn_tco38: string;
   attribute syn_tco38 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[8] = 3.908";
   attribute syn_tco39: string;
   attribute syn_tco39 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[9] = 3.932";
   attribute syn_tco40: string;
   attribute syn_tco40 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_READYOUT = 3.615";
   attribute syn_tco41: string;
   attribute syn_tco41 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RESP = 3.751";
   attribute syn_tco42: string;
   attribute syn_tco42 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[0] = 3.660";
   attribute syn_tco43: string;
   attribute syn_tco43 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[10] = 3.949";
   attribute syn_tco44: string;
   attribute syn_tco44 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[11] = 3.596";
   attribute syn_tco45: string;
   attribute syn_tco45 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[12] = 3.677";
   attribute syn_tco46: string;
   attribute syn_tco46 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[13] = 3.647";
   attribute syn_tco47: string;
   attribute syn_tco47 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[14] = 3.652";
   attribute syn_tco48: string;
   attribute syn_tco48 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[15] = 3.580";
   attribute syn_tco49: string;
   attribute syn_tco49 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[16] = 3.611";
   attribute syn_tco50: string;
   attribute syn_tco50 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[17] = 3.697";
   attribute syn_tco51: string;
   attribute syn_tco51 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[18] = 3.696";
   attribute syn_tco52: string;
   attribute syn_tco52 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[19] = 3.893";
   attribute syn_tco53: string;
   attribute syn_tco53 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[1] = 3.597";
   attribute syn_tco54: string;
   attribute syn_tco54 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[20] = 3.631";
   attribute syn_tco55: string;
   attribute syn_tco55 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[21] = 3.748";
   attribute syn_tco56: string;
   attribute syn_tco56 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[22] = 3.686";
   attribute syn_tco57: string;
   attribute syn_tco57 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[23] = 3.709";
   attribute syn_tco58: string;
   attribute syn_tco58 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[24] = 3.730";
   attribute syn_tco59: string;
   attribute syn_tco59 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[25] = 3.555";
   attribute syn_tco60: string;
   attribute syn_tco60 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[26] = 3.854";
   attribute syn_tco61: string;
   attribute syn_tco61 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[27] = 3.732";
   attribute syn_tco62: string;
   attribute syn_tco62 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[28] = 4.096";
   attribute syn_tco63: string;
   attribute syn_tco63 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[29] = 3.532";
   attribute syn_tco64: string;
   attribute syn_tco64 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[2] = 3.576";
   attribute syn_tco65: string;
   attribute syn_tco65 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[30] = 3.519";
   attribute syn_tco66: string;
   attribute syn_tco66 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[31] = 3.889";
   attribute syn_tco67: string;
   attribute syn_tco67 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[3] = 3.576";
   attribute syn_tco68: string;
   attribute syn_tco68 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[4] = 3.560";
   attribute syn_tco69: string;
   attribute syn_tco69 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[5] = 3.657";
   attribute syn_tco70: string;
   attribute syn_tco70 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[6] = 3.746";
   attribute syn_tco71: string;
   attribute syn_tco71 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[7] = 3.593";
   attribute syn_tco72: string;
   attribute syn_tco72 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[8] = 3.945";
   attribute syn_tco73: string;
   attribute syn_tco73 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[9] = 3.735";
   attribute syn_tco74: string;
   attribute syn_tco74 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ENABLE = 3.736";
   attribute syn_tco75: string;
   attribute syn_tco75 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SEL = 3.488";
   attribute syn_tco76: string;
   attribute syn_tco76 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[0] = 3.648";
   attribute syn_tco77: string;
   attribute syn_tco77 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[10] = 3.504";
   attribute syn_tco78: string;
   attribute syn_tco78 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[11] = 3.726";
   attribute syn_tco79: string;
   attribute syn_tco79 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[12] = 3.725";
   attribute syn_tco80: string;
   attribute syn_tco80 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[13] = 3.782";
   attribute syn_tco81: string;
   attribute syn_tco81 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[14] = 3.722";
   attribute syn_tco82: string;
   attribute syn_tco82 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[15] = 3.787";
   attribute syn_tco83: string;
   attribute syn_tco83 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[16] = 3.624";
   attribute syn_tco84: string;
   attribute syn_tco84 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[17] = 3.878";
   attribute syn_tco85: string;
   attribute syn_tco85 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[18] = 3.653";
   attribute syn_tco86: string;
   attribute syn_tco86 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[19] = 3.811";
   attribute syn_tco87: string;
   attribute syn_tco87 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[1] = 3.743";
   attribute syn_tco88: string;
   attribute syn_tco88 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[20] = 3.672";
   attribute syn_tco89: string;
   attribute syn_tco89 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[21] = 3.625";
   attribute syn_tco90: string;
   attribute syn_tco90 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[22] = 3.639";
   attribute syn_tco91: string;
   attribute syn_tco91 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[23] = 3.628";
   attribute syn_tco92: string;
   attribute syn_tco92 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[24] = 3.784";
   attribute syn_tco93: string;
   attribute syn_tco93 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[25] = 3.361";
   attribute syn_tco94: string;
   attribute syn_tco94 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[26] = 3.699";
   attribute syn_tco95: string;
   attribute syn_tco95 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[27] = 3.382";
   attribute syn_tco96: string;
   attribute syn_tco96 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[28] = 3.753";
   attribute syn_tco97: string;
   attribute syn_tco97 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[29] = 3.423";
   attribute syn_tco98: string;
   attribute syn_tco98 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[2] = 3.769";
   attribute syn_tco99: string;
   attribute syn_tco99 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[30] = 3.735";
   attribute syn_tco100: string;
   attribute syn_tco100 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[31] = 3.364";
   attribute syn_tco101: string;
   attribute syn_tco101 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[3] = 3.838";
   attribute syn_tco102: string;
   attribute syn_tco102 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[4] = 3.566";
   attribute syn_tco103: string;
   attribute syn_tco103 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[5] = 3.656";
   attribute syn_tco104: string;
   attribute syn_tco104 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[6] = 3.667";
   attribute syn_tco105: string;
   attribute syn_tco105 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[7] = 3.881";
   attribute syn_tco106: string;
   attribute syn_tco106 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[8] = 3.612";
   attribute syn_tco107: string;
   attribute syn_tco107 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[9] = 3.648";
   attribute syn_tco108: string;
   attribute syn_tco108 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WRITE = 3.682";
   attribute syn_tco109: string;
   attribute syn_tco109 of DEF_ARCH : architecture is " CLK_BASE->H2FCALIB = 3.640";
   attribute syn_tco110: string;
   attribute syn_tco110 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_MGPIO31B_H2F_B = 3.188";
   attribute syn_tco111: string;
   attribute syn_tco111 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_USBC_DATA1_MGPIO31B_OE = 3.985";
   attribute syn_tco112: string;
   attribute syn_tco112 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_A = 3.182";
   attribute syn_tco113: string;
   attribute syn_tco113 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_B = 3.192";
   attribute syn_tco114: string;
   attribute syn_tco114 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_USBC_DATA0_MGPIO30B_OE = 3.772";
   attribute syn_tco115: string;
   attribute syn_tco115 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_MGPIO1A_H2F_B = 3.346";
   attribute syn_tco116: string;
   attribute syn_tco116 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_USBA_DATA4_MGPIO1A_OE = 3.478";
   attribute syn_tco117: string;
   attribute syn_tco117 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_A = 3.284";
   attribute syn_tco118: string;
   attribute syn_tco118 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_B = 3.436";
   attribute syn_tco119: string;
   attribute syn_tco119 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_USBA_DATA3_MGPIO0A_OE = 3.212";
   attribute syn_tco120: string;
   attribute syn_tco120 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_A = 3.383";
   attribute syn_tco121: string;
   attribute syn_tco121 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_B = 3.249";
   attribute syn_tco122: string;
   attribute syn_tco122 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_A = 3.254";
   attribute syn_tco123: string;
   attribute syn_tco123 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_B = 3.219";
   attribute syn_tco124: string;
   attribute syn_tco124 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_A = 3.239";
   attribute syn_tco125: string;
   attribute syn_tco125 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_B = 3.270";
   attribute syn_tco126: string;
   attribute syn_tco126 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_A = 3.307";
   attribute syn_tco127: string;
   attribute syn_tco127 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_B = 3.259";
   attribute syn_tco128: string;
   attribute syn_tco128 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT = 3.335";
   attribute syn_tco129: string;
   attribute syn_tco129 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_A = 3.320";
   attribute syn_tco130: string;
   attribute syn_tco130 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_B = 3.255";
   attribute syn_tco131: string;
   attribute syn_tco131 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_A = 3.313";
   attribute syn_tco132: string;
   attribute syn_tco132 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_B = 3.330";
   attribute syn_tco133: string;
   attribute syn_tco133 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT = 3.332";
   attribute syn_tco134: string;
   attribute syn_tco134 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_A = 3.253";
   attribute syn_tco135: string;
   attribute syn_tco135 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_B = 3.152";
   attribute syn_tco136: string;
   attribute syn_tco136 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_A = 3.246";
   attribute syn_tco137: string;
   attribute syn_tco137 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_B = 3.213";
   attribute syn_tco138: string;
   attribute syn_tco138 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OE = 3.789";
   attribute syn_tco139: string;
   attribute syn_tco139 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OUT = 3.182";
   attribute syn_tco140: string;
   attribute syn_tco140 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_A = 3.878";
   attribute syn_tco141: string;
   attribute syn_tco141 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_B = 3.928";
   attribute syn_tco142: string;
   attribute syn_tco142 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OE = 3.813";
   attribute syn_tco143: string;
   attribute syn_tco143 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OUT = 3.494";
   attribute syn_tco144: string;
   attribute syn_tco144 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_H2F_A = 3.262";
   attribute syn_tco145: string;
   attribute syn_tco145 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_A = 3.252";
   attribute syn_tco146: string;
   attribute syn_tco146 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_B = 3.279";
   attribute syn_tco147: string;
   attribute syn_tco147 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_A = 3.206";
   attribute syn_tco148: string;
   attribute syn_tco148 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_B = 3.113";
   attribute syn_tco149: string;
   attribute syn_tco149 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_A = 3.342";
   attribute syn_tco150: string;
   attribute syn_tco150 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_B = 3.278";
   attribute syn_tco151: string;
   attribute syn_tco151 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OE = 3.543";
   attribute syn_tco152: string;
   attribute syn_tco152 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT = 3.221";
   attribute syn_tco153: string;
   attribute syn_tco153 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_A = 3.206";
   attribute syn_tco154: string;
   attribute syn_tco154 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_B = 3.228";
   attribute syn_tco155: string;
   attribute syn_tco155 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OE = 3.798";
   attribute syn_tco156: string;
   attribute syn_tco156 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT = 3.509";
   attribute syn_tco157: string;
   attribute syn_tco157 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE = 1.207";
   attribute syn_tco158: string;
   attribute syn_tco158 of DEF_ARCH : architecture is " CLK_BASE->RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE = 1.588";
   attribute syn_tco159: string;
   attribute syn_tco159 of DEF_ARCH : architecture is " CLK_BASE->RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE = 1.189";
   attribute syn_tco160: string;
   attribute syn_tco160 of DEF_ARCH : architecture is " CLK_BASE->RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE = 1.213";
   attribute syn_tco161: string;
   attribute syn_tco161 of DEF_ARCH : architecture is " CLK_BASE->RGMII_RXD3_USBB_DATA4_OE = 1.246";
   attribute syn_tco162: string;
   attribute syn_tco162 of DEF_ARCH : architecture is " CLK_BASE->RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE = 1.257";
   attribute syn_tco163: string;
   attribute syn_tco163 of DEF_ARCH : architecture is " CLK_BASE->RGMII_TXD1_RMII_TXD1_USBB_STP_OUT = 4.390";
   attribute syn_tco164: string;
   attribute syn_tco164 of DEF_ARCH : architecture is " CLK_BASE->RGMII_TXD2_USBB_DATA5_OE = 1.128";
   attribute syn_tco165: string;
   attribute syn_tco165 of DEF_ARCH : architecture is " CLK_BASE->RGMII_TXD3_USBB_DATA6_OE = 0.841";
   attribute syn_tco166: string;
   attribute syn_tco166 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_A = 3.181";
   attribute syn_tco167: string;
   attribute syn_tco167 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_B = 3.251";
   attribute syn_tco168: string;
   attribute syn_tco168 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_A = 3.287";
   attribute syn_tco169: string;
   attribute syn_tco169 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_B = 3.353";
   attribute syn_tco170: string;
   attribute syn_tco170 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OE = 5.073";
   attribute syn_tco171: string;
   attribute syn_tco171 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OUT = 5.638";
   attribute syn_tco172: string;
   attribute syn_tco172 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_A = 3.240";
   attribute syn_tco173: string;
   attribute syn_tco173 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_B = 3.270";
   attribute syn_tco174: string;
   attribute syn_tco174 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_A = 3.262";
   attribute syn_tco175: string;
   attribute syn_tco175 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_B = 3.303";
   attribute syn_tco176: string;
   attribute syn_tco176 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_A = 3.237";
   attribute syn_tco177: string;
   attribute syn_tco177 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_B = 3.267";
   attribute syn_tco178: string;
   attribute syn_tco178 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_A = 3.187";
   attribute syn_tco179: string;
   attribute syn_tco179 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_B = 3.112";
   attribute syn_tco180: string;
   attribute syn_tco180 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS4_MGPIO19A_H2F_A = 3.215";
   attribute syn_tco181: string;
   attribute syn_tco181 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS5_MGPIO20A_H2F_A = 3.345";
   attribute syn_tco182: string;
   attribute syn_tco182 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS6_MGPIO21A_H2F_A = 3.385";
   attribute syn_tco183: string;
   attribute syn_tco183 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS7_MGPIO22A_H2F_A = 3.320";
   attribute syn_tco184: string;
   attribute syn_tco184 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_A = 3.253";
   attribute syn_tco185: string;
   attribute syn_tco185 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_B = 3.201";
   attribute syn_tco186: string;
   attribute syn_tco186 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_A = 3.174";
   attribute syn_tco187: string;
   attribute syn_tco187 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_B = 3.251";
   attribute syn_tco188: string;
   attribute syn_tco188 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OE = 5.581";
   attribute syn_tco189: string;
   attribute syn_tco189 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OUT = 6.229";
   attribute syn_tco190: string;
   attribute syn_tco190 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_A = 3.204";
   attribute syn_tco191: string;
   attribute syn_tco191 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_B = 3.183";
   attribute syn_tco192: string;
   attribute syn_tco192 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_A = 3.223";
   attribute syn_tco193: string;
   attribute syn_tco193 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_B = 3.291";
   attribute syn_tco194: string;
   attribute syn_tco194 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_A = 3.345";
   attribute syn_tco195: string;
   attribute syn_tco195 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_B = 3.261";
   attribute syn_tco196: string;
   attribute syn_tco196 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_A = 3.270";
   attribute syn_tco197: string;
   attribute syn_tco197 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_B = 3.378";
   attribute syn_tco198: string;
   attribute syn_tco198 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS4_MGPIO17A_H2F_A = 3.245";
   attribute syn_tco199: string;
   attribute syn_tco199 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS5_MGPIO18A_H2F_A = 3.282";
   attribute syn_tco200: string;
   attribute syn_tco200 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS6_MGPIO23A_H2F_A = 3.253";
   attribute syn_tco201: string;
   attribute syn_tco201 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS7_MGPIO24A_H2F_A = 3.232";
   attribute black_box_pad_pin : string;
   attribute black_box_pad_pin of DEF_ARCH : architecture is "";

begin

end DEF_ARCH;
